module codememory_sort(c1,readselect,writeselect,inp,outp,clk,reset);
	input wire c1,clk,reset;input wire[5:0]readselect,writeselect;
	input wire [15:0]inp;
	output wire [15:0]outp;
	reg [15:0] c [0:63];
	
	
	always @(posedge clk , posedge reset) begin
		if (reset) begin
			c[0]  = 16'b0000000000000000;
			c[1]  = 16'b1110_00_00_00011110;//jump to 32
			c[2]  = 16'b0000000000000000;
			c[3]  = 16'b0000000000000000;
			c[4]  = 16'b0000000000000000;
			c[5]  = 16'b0000000000000000;
			c[6]  = 16'b0000000000000000;
			c[7]  = 16'b0000000000000000;
			c[8]  = 16'b0000000000000000;
			c[9]  = 16'b0000000000000000;
			c[10] = 16'b0000000000000000;
			c[11] = 16'b0000000000000000;
			c[12] = 16'b0000000000000000;
			c[13] = 16'b0000000000000000;
			c[14] = 16'b0000000000000000;
			c[15] = 16'b0000000000000000;
			c[16] = 16'b0000000000000000;
			c[17] = 16'b0000000000000000;
			c[18] = 16'b0000000000000000;
			c[19] = 16'b0000000000000000;
			c[20] = 16'b0000000000000000;
			c[21] = 16'b0000000000000000;
			c[22] = 16'b0000000000000000;
			c[23] = 16'b0000000000000000;
			c[24] = 16'b0000000000000000;
			c[25] = 16'b0000000000000000;
			c[26] = 16'b0000000000000000;
			c[27] = 16'b0000000000000000;
			c[28] = 16'b0000000000000000;
			c[29] = 16'b0000000000000000;
			c[30] = 16'b0000000000000000;
			c[31] = 16'b0000000000000000;
			c[32] = 16'b0011000000000000; // LOADI  A  ,  0
			c[33] = 16'b1000110000001000; // Outer:  LOAD   D  ,   [  last  ]
			c[34] = 16'b0011010000000000; // LOADI  B  ,  0
			c[35] = 16'b1101001100000000; // CMP    A  ,  D
			c[36] = 16'b1111001100001110; // BRGE   End
			c[37] = 16'b1000110000001000; // Inner:  LOAD   D  ,   [  last  ]
			c[38] = 16'b0110110000000000; // SUB    D  ,  A
			c[39] = 16'b1101011100000000; // CMP    B  ,  D
			c[40] = 16'b1111001100001000; // BRGE   Iinc
			c[41] = 16'b1001100100000000; // If:     LOADF  C  ,   [  array  +  B  ]
			c[42] = 16'b1001110100000001; //         LOADF  D  ,   [  array  +  B  +  1  ]
			c[43] = 16'b1101111000000000; //         CMP    D  ,  C
			c[44] = 16'b1111001100000010; //         BRGE   Jinc
			c[45] = 16'b1011110100000000; // Swap:   STOREF  [  array  +  B  ]   ,  D
			c[46] = 16'b1011100100000001; //         STOREF  [  array  +  B  +  1  ]   ,  C
			c[47] = 16'b0101010000000001; // Jinc:   ADDI   B  ,  1
			c[48]  = 16'b1110000011110100; // JUMP   Inner
			c[49]  = 16'b0101000000000001; // Iinc:   ADDI   A  ,  1
			c[50]  = 16'b1110000011101110; // JUMP   Outer
			c[51]  = 16'b0000000000000000; // End:    NOOP
			c[52]  = 16'b0000000000000000;
			c[53]  = 16'b0000000000000000;
			c[54]  = 16'b0000000000000000;
			c[55]  = 16'b0000000000000000;
			c[56]  = 16'b0000000000000000;
			c[57]  = 16'b0000000000000000;
			c[58]  = 16'b0000000000000000;
			c[59]  = 16'b0000000000000000;
			c[60]  = 16'b0000000000000000;
			c[61]  = 16'b0000000000000000;
			c[62]  = 16'b0000000000000000;
			c[63]  = 16'b0000000000000000;
		end
		else begin
			if(c1==1'b1)
				c[writeselect] <= inp;
		end
	end
	
	assign outp = c[readselect];
	
endmodule 